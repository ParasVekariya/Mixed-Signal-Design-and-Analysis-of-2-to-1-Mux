* /home/paras.vekariya/eSim-Workspace/mixed/mixed.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri 07 Oct 2022 08:11:13 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ parasvekariya_2in1mux		
v3  select GND pulse		
v2  D1 GND pulse		
v1  D0 GND pulse		
U3  select plot_v1		
U2  D1 plot_v1		
U1  D0 plot_v1		
U5  D0 D1 select Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ adc_bridge_3		
U6  Net-_U4-Pad4_ Net-_SC1-Pad1_ dac_bridge_1		
SC1  Net-_SC1-Pad1_ Y_out Net-_SC1-Pad1_ sky130_fd_pr__res_generic_pd		
SC2  Y_out GND sky130_fd_pr__cap_mim_m3_1		
U7  Y_out plot_v1		
scmode1  SKY130mode		

.end
